package fsm_pkg;
	typedef enum int unsigned {IDLE,
							   START,
                               VIEW,
                               NVIEW,
							   XXX} state_e;
endpackage: fsm_pkg